class i2c_scoreboard_freq extends uvm_scoreboard;
  `uvm_component_utils(i2c_scoreboard_freq)

endclass : i2c_scoreboard_freq
